component traffic_light.CDiagnosticsMessage

endpoints {
    dmessage : traffic_light.IDiagnosticsMessage
}