component traffic_light.DiagnosticsMessage

endpoints {
    dmessage : traffic_light.DiagnosticsMessage
}